module INV (A, F);
	assign F = ~A;
endmodule