module top;
	initial begin
	 $display ( "Hello World!" );
	end
endmodule
