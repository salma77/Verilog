module INV (A, F);
	input A;
	output F;
	assign F = ~A;
endmodule