module FULLADD ();
//How will it take a vector?!
endmodule
